picorv32/picorv32.v