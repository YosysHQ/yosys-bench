picorv32/scripts/vivado/synth_area_top.v