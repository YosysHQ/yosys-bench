picorv32/picosoc/picosoc.v