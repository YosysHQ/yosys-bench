picorv32/picosoc/simpleuart.v