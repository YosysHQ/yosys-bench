picorv32/picosoc/spimemio.v